module TreeLUT(input wire [53:0] i, output wire [20:0] o);


wire [50:0] binary_features;

assign binary_features[0] = (i[0:0] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[1] = (i[1:1] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[2] = (i[2:2] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[3] = (i[3:3] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[4] = (i[4:4] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[5] = (i[5:5] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[6] = (i[6:6] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[7] = (i[7:7] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[8] = (i[8:8] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[9] = (i[9:9] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[10] = (i[10:10] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[11] = (i[11:11] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[12] = (i[12:12] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[13] = (i[13:13] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[14] = (i[14:14] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[15] = (i[15:15] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[16] = (i[16:16] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[17] = (i[19:19] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[18] = (i[20:20] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[19] = (i[21:21] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[20] = (i[22:22] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[21] = (i[23:23] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[22] = (i[24:24] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[23] = (i[26:26] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[24] = (i[27:27] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[25] = (i[28:28] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[26] = (i[29:29] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[27] = (i[30:30] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[28] = (i[31:31] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[29] = (i[32:32] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[30] = (i[33:33] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[31] = (i[34:34] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[32] = (i[35:35] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[33] = (i[36:36] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[34] = (i[37:37] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[35] = (i[38:38] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[36] = (i[39:39] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[37] = (i[40:40] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[38] = (i[41:41] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[39] = (i[42:42] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[40] = (i[43:43] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[41] = (i[44:44] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[42] = (i[45:45] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[43] = (i[46:46] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[44] = (i[47:47] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[45] = (i[48:48] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[46] = (i[49:49] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[47] = (i[50:50] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[48] = (i[51:51] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[49] = (i[52:52] < (1'd1))? 1'b1 : 1'b0;
assign binary_features[50] = (i[53:53] < (1'd1))? 1'b1 : 1'b0;


wire [48:0] trees_output;

class0_tree0 class0_tree0_inst(.i(binary_features), .o(trees_output[0:0]));
class0_tree1 class0_tree1_inst(.i(binary_features), .o(trees_output[1:1]));
class0_tree2 class0_tree2_inst(.i(binary_features), .o(trees_output[2:2]));
class0_tree3 class0_tree3_inst(.i(binary_features), .o(trees_output[3:3]));
class0_tree4 class0_tree4_inst(.i(binary_features), .o(trees_output[4:4]));
class0_tree5 class0_tree5_inst(.i(binary_features), .o(trees_output[5:5]));
class0_tree6 class0_tree6_inst(.i(binary_features), .o(trees_output[6:6]));
class1_tree0 class1_tree0_inst(.i(binary_features), .o(trees_output[7:7]));
class1_tree1 class1_tree1_inst(.i(binary_features), .o(trees_output[8:8]));
class1_tree2 class1_tree2_inst(.i(binary_features), .o(trees_output[9:9]));
class1_tree3 class1_tree3_inst(.i(binary_features), .o(trees_output[10:10]));
class1_tree4 class1_tree4_inst(.i(binary_features), .o(trees_output[11:11]));
class1_tree5 class1_tree5_inst(.i(binary_features), .o(trees_output[12:12]));
class1_tree6 class1_tree6_inst(.i(binary_features), .o(trees_output[13:13]));
class2_tree0 class2_tree0_inst(.i(binary_features), .o(trees_output[14:14]));
class2_tree1 class2_tree1_inst(.i(binary_features), .o(trees_output[15:15]));
class2_tree2 class2_tree2_inst(.i(binary_features), .o(trees_output[16:16]));
class2_tree3 class2_tree3_inst(.i(binary_features), .o(trees_output[17:17]));
class2_tree4 class2_tree4_inst(.i(binary_features), .o(trees_output[18:18]));
class2_tree5 class2_tree5_inst(.i(binary_features), .o(trees_output[19:19]));
class2_tree6 class2_tree6_inst(.i(binary_features), .o(trees_output[20:20]));
class3_tree0 class3_tree0_inst(.i(binary_features), .o(trees_output[21:21]));
class3_tree1 class3_tree1_inst(.i(binary_features), .o(trees_output[22:22]));
class3_tree2 class3_tree2_inst(.i(binary_features), .o(trees_output[23:23]));
class3_tree3 class3_tree3_inst(.i(binary_features), .o(trees_output[24:24]));
class3_tree4 class3_tree4_inst(.i(binary_features), .o(trees_output[25:25]));
class3_tree5 class3_tree5_inst(.i(binary_features), .o(trees_output[26:26]));
class3_tree6 class3_tree6_inst(.i(binary_features), .o(trees_output[27:27]));
class4_tree0 class4_tree0_inst(.i(binary_features), .o(trees_output[28:28]));
class4_tree1 class4_tree1_inst(.i(binary_features), .o(trees_output[29:29]));
class4_tree2 class4_tree2_inst(.i(binary_features), .o(trees_output[30:30]));
class4_tree3 class4_tree3_inst(.i(binary_features), .o(trees_output[31:31]));
class4_tree4 class4_tree4_inst(.i(binary_features), .o(trees_output[32:32]));
class4_tree5 class4_tree5_inst(.i(binary_features), .o(trees_output[33:33]));
class4_tree6 class4_tree6_inst(.i(binary_features), .o(trees_output[34:34]));
class5_tree0 class5_tree0_inst(.i(binary_features), .o(trees_output[35:35]));
class5_tree1 class5_tree1_inst(.i(binary_features), .o(trees_output[36:36]));
class5_tree2 class5_tree2_inst(.i(binary_features), .o(trees_output[37:37]));
class5_tree3 class5_tree3_inst(.i(binary_features), .o(trees_output[38:38]));
class5_tree4 class5_tree4_inst(.i(binary_features), .o(trees_output[39:39]));
class5_tree5 class5_tree5_inst(.i(binary_features), .o(trees_output[40:40]));
class5_tree6 class5_tree6_inst(.i(binary_features), .o(trees_output[41:41]));
class6_tree0 class6_tree0_inst(.i(binary_features), .o(trees_output[42:42]));
class6_tree1 class6_tree1_inst(.i(binary_features), .o(trees_output[43:43]));
class6_tree2 class6_tree2_inst(.i(binary_features), .o(trees_output[44:44]));
class6_tree3 class6_tree3_inst(.i(binary_features), .o(trees_output[45:45]));
class6_tree4 class6_tree4_inst(.i(binary_features), .o(trees_output[46:46]));
class6_tree5 class6_tree5_inst(.i(binary_features), .o(trees_output[47:47]));
class6_tree6 class6_tree6_inst(.i(binary_features), .o(trees_output[48:48]));

class0_adder class0_adder_inst(.i(trees_output[6:0]), .o(o[2:0]));
class1_adder class1_adder_inst(.i(trees_output[13:7]), .o(o[5:3]));
class2_adder class2_adder_inst(.i(trees_output[20:14]), .o(o[8:6]));
class3_adder class3_adder_inst(.i(trees_output[27:21]), .o(o[11:9]));
class4_adder class4_adder_inst(.i(trees_output[34:28]), .o(o[14:12]));
class5_adder class5_adder_inst(.i(trees_output[41:35]), .o(o[17:15]));
class6_adder class6_adder_inst(.i(trees_output[48:42]), .o(o[20:18]));

endmodule
