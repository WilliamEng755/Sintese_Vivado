module class6_tree6(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_36;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_44;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_52;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_57;
wire [0:0] new_59;
wire [0:0] new_60;
wire [0:0] new_61;
wire [0:0] new_62;
wire [0:0] new_63;
wire [0:0] new_64;
assign new_64 = i[4] ? 0 : 0;
assign new_63 = i[2] ? 0 : 0;
assign new_62 = i[2] ? 0 : 0;
assign new_61 = i[2] ? 0 : 0;
assign new_60 = i[5] ? 0 : 0;
assign new_59 = i[5] ? 0 : 0;
assign new_57 = i[0] ? 0 : 0;
assign new_55 = i[9] ? 0 : 0;
assign new_54 = i[0] ? 0 : 0;
assign new_53 = i[8] ? 0 : 0;
assign new_52 = i[5] ? 0 : 0;
assign new_51 = i[48] ? 0 : 0;
assign new_50 = i[4] ? 0 : 0;
assign new_48 = i[9] ? 0 : 0;
assign new_47 = i[0] ? 0 : 0;
assign new_46 = i[4] ? 0 : 0;
assign new_45 = i[3] ? 0 : 0;
assign new_44 = i[3] ? 0 : 0;
assign new_43 = i[3] ? 0 : 0;
assign new_42 = i[3] ? 0 : 0;
assign new_41 = i[4] ? 0 : 0;
assign new_39 = i[1] ? 0 : 0;
assign new_38 = i[8] ? 0 : 0;
assign new_36 = i[8] ? 0 : 0;
assign new_35 = i[1] ? 0 : 0;
assign new_34 = i[4] ? 0 : 0;
assign new_33 = i[49] ? 0 : 0;
assign new_32 = i[8] ? new_63 : new_64;
assign new_31 = i[5] ? new_61 : new_62;
assign new_30 = i[3] ? new_59 : new_60;
assign new_29 = i[2] ? new_57 : 0;
assign new_28 = i[4] ? new_55 : 0;
assign new_27 = i[3] ? new_53 : new_54;
assign new_26 = i[3] ? new_51 : new_52;
assign new_25 = i[6] ? 0 : new_50;
assign new_24 = i[4] ? new_47 : new_48;
assign new_23 = i[5] ? new_45 : new_46;
assign new_22 = i[8] ? new_43 : new_44;
assign new_21 = i[8] ? new_41 : new_42;
assign new_20 = i[2] ? new_39 : 0;
assign new_19 = i[6] ? 0 : new_38;
assign new_18 = i[48] ? new_35 : new_36;
assign new_17 = i[43] ? new_33 : new_34;
assign new_16 = i[1] ? new_31 : new_32;
assign new_15 = i[9] ? new_29 : new_30;
assign new_14 = i[48] ? new_27 : new_28;
assign new_13 = i[0] ? new_25 : new_26;
assign new_12 = i[8] ? new_23 : new_24;
assign new_11 = i[5] ? new_21 : new_22;
assign new_10 = i[49] ? new_19 : new_20;
assign new_9 = i[42] ? new_17 : new_18;
assign new_8 = i[6] ? new_15 : new_16;
assign new_7 = i[2] ? new_13 : new_14;
assign new_6 = i[49] ? new_11 : new_12;
assign new_5 = i[47] ? new_9 : new_10;
assign new_4 = i[10] ? new_7 : new_8;
assign new_3 = i[45] ? new_5 : new_6;
assign new_1 = i[46] ? new_3 : new_4;
assign o = i[50] ? new_1 : 0;


endmodule
