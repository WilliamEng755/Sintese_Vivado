module class1_tree4(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_36;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_49;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_52;
wire [0:0] new_54;
wire [0:0] new_57;
wire [0:0] new_59;
wire [0:0] new_60;
wire [0:0] new_61;
wire [0:0] new_62;
wire [0:0] new_63;
wire [0:0] new_64;
wire [0:0] new_65;
wire [0:0] new_67;
wire [0:0] new_69;
wire [0:0] new_71;
wire [0:0] new_73;
wire [0:0] new_74;
wire [0:0] new_75;
wire [0:0] new_77;
wire [0:0] new_78;
wire [0:0] new_79;
wire [0:0] new_81;
wire [0:0] new_82;
wire [0:0] new_83;
wire [0:0] new_84;
wire [0:0] new_85;
wire [0:0] new_86;
wire [0:0] new_87;
wire [0:0] new_89;
wire [0:0] new_90;
wire [0:0] new_92;
assign new_92 = i[9] ? 0 : 0;
assign new_90 = i[0] ? 0 : 0;
assign new_89 = i[1] ? 0 : 0;
assign new_87 = i[0] ? 0 : 0;
assign new_86 = i[4] ? 0 : 0;
assign new_85 = i[3] ? 0 : 0;
assign new_84 = i[0] ? 0 : 0;
assign new_83 = i[0] ? 0 : 0;
assign new_82 = i[1] ? 0 : 0;
assign new_81 = i[5] ? 0 : 0;
assign new_79 = i[5] ? 0 : 0;
assign new_78 = i[3] ? 0 : 0;
assign new_77 = i[4] ? 0 : 0;
assign new_75 = i[8] ? 0 : 0;
assign new_74 = i[1] ? 0 : 0;
assign new_73 = i[4] ? 0 : 0;
assign new_71 = i[9] ? 0 : 0;
assign new_69 = i[9] ? 0 : 0;
assign new_67 = i[3] ? 0 : 0;
assign new_65 = i[5] ? 0 : 0;
assign new_64 = i[0] ? 0 : 0;
assign new_63 = i[4] ? 0 : 0;
assign new_62 = i[1] ? 0 : 0;
assign new_61 = i[4] ? 0 : 0;
assign new_60 = i[1] ? 0 : 0;
assign new_59 = i[0] ? 0 : 0;
assign new_57 = i[41] ? 0 : 0;
assign new_54 = i[1] ? 0 : new_92;
assign new_52 = i[4] ? new_89 : new_90;
assign new_51 = i[3] ? new_87 : 0;
assign new_50 = i[5] ? new_85 : new_86;
assign new_49 = i[3] ? new_83 : new_84;
assign new_48 = i[3] ? new_81 : new_82;
assign new_47 = i[1] ? new_79 : 0;
assign new_46 = i[9] ? new_77 : new_78;
assign new_43 = i[1] ? new_75 : 0;
assign new_42 = i[8] ? new_73 : new_74;
assign new_41 = i[8] ? new_71 : 0;
assign new_39 = i[5] ? new_69 : 0;
assign new_38 = i[5] ? new_67 : 0;
assign new_36 = i[3] ? new_65 : 0;
assign new_34 = i[1] ? new_63 : new_64;
assign new_33 = i[0] ? new_61 : new_62;
assign new_32 = i[48] ? new_59 : new_60;
assign new_31 = i[11] ? new_57 : 0;
assign new_30 = i[9] ? 0 : 0;
assign new_29 = i[8] ? 0 : new_54;
assign new_26 = i[8] ? new_51 : new_52;
assign new_25 = i[1] ? new_49 : new_50;
assign new_24 = i[8] ? new_47 : new_48;
assign new_23 = i[8] ? 0 : new_46;
assign new_22 = i[5] ? new_43 : 0;
assign new_21 = i[5] ? new_41 : new_42;
assign new_20 = i[1] ? new_39 : 0;
assign new_19 = i[8] ? 0 : new_38;
assign new_18 = i[48] ? 0 : new_36;
assign new_16 = i[8] ? new_33 : new_34;
assign new_15 = i[45] ? new_31 : new_32;
assign new_14 = i[3] ? new_29 : new_30;
assign new_13 = i[1] ? 0 : 0;
assign new_12 = i[9] ? new_25 : new_26;
assign new_11 = i[0] ? new_23 : new_24;
assign new_10 = i[3] ? new_21 : new_22;
assign new_9 = i[4] ? new_19 : new_20;
assign new_8 = i[1] ? 0 : new_18;
assign new_7 = i[33] ? new_15 : new_16;
assign new_6 = i[4] ? new_13 : new_14;
assign new_5 = i[10] ? new_11 : new_12;
assign new_4 = i[0] ? new_9 : new_10;
assign new_3 = i[42] ? new_7 : new_8;
assign new_2 = i[48] ? new_5 : new_6;
assign new_1 = i[17] ? new_3 : new_4;
assign o = i[26] ? new_1 : new_2;


endmodule
