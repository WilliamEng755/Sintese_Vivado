module class0_tree2(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_37;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_50;
wire [0:0] new_52;
assign new_52 = i[8] ? 0 : 0;
assign new_50 = i[8] ? 0 : 0;
assign new_48 = i[4] ? 0 : 0;
assign new_47 = i[26] ? 0 : 0;
assign new_43 = i[14] ? 0 : 0;
assign new_42 = i[5] ? 0 : 0;
assign new_41 = i[6] ? 0 : 0;
assign new_40 = i[5] ? 0 : 0;
assign new_39 = i[3] ? 0 : 0;
assign new_38 = i[3] ? 0 : 0;
assign new_37 = i[0] ? 0 : 0;
assign new_35 = i[3] ? 0 : 0;
assign new_34 = i[3] ? 0 : 0;
assign new_33 = i[48] ? 0 : 0;
assign new_32 = i[8] ? 0 : 0;
assign new_31 = i[21] ? 0 : 0;
assign new_30 = i[4] ? 0 : new_52;
assign new_29 = i[4] ? 0 : new_50;
assign new_27 = i[39] ? new_47 : new_48;
assign new_26 = i[4] ? 0 : 0;
assign new_25 = i[41] ? new_43 : 0;
assign new_24 = i[4] ? new_41 : new_42;
assign new_23 = i[4] ? new_39 : new_40;
assign new_22 = i[9] ? new_37 : new_38;
assign new_21 = i[5] ? new_35 : 0;
assign new_18 = i[8] ? new_33 : new_34;
assign new_17 = i[19] ? new_31 : new_32;
assign new_16 = i[0] ? new_29 : new_30;
assign new_15 = i[38] ? new_27 : 0;
assign new_13 = i[13] ? new_25 : new_26;
assign new_12 = i[0] ? new_23 : new_24;
assign new_11 = i[4] ? new_21 : new_22;
assign new_10 = i[10] ? 0 : 0;
assign new_9 = i[30] ? new_17 : new_18;
assign new_8 = i[40] ? new_15 : new_16;
assign new_7 = i[33] ? new_13 : 0;
assign new_6 = i[8] ? new_11 : new_12;
assign new_5 = i[25] ? new_9 : new_10;
assign new_4 = i[48] ? new_7 : new_8;
assign new_3 = i[18] ? new_5 : new_6;
assign new_1 = i[1] ? new_3 : new_4;
assign o = i[50] ? new_1 : 0;


endmodule
