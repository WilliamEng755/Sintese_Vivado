module class6_tree4(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_36;
wire [0:0] new_37;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_44;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_49;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_52;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_57;
wire [0:0] new_59;
wire [0:0] new_60;
wire [0:0] new_61;
wire [0:0] new_63;
wire [0:0] new_65;
wire [0:0] new_66;
wire [0:0] new_67;
wire [0:0] new_68;
wire [0:0] new_69;
wire [0:0] new_70;
wire [0:0] new_71;
wire [0:0] new_72;
wire [0:0] new_73;
wire [0:0] new_74;
wire [0:0] new_75;
wire [0:0] new_76;
wire [0:0] new_77;
wire [0:0] new_79;
wire [0:0] new_80;
wire [0:0] new_81;
wire [0:0] new_82;
wire [0:0] new_84;
wire [0:0] new_85;
wire [0:0] new_87;
wire [0:0] new_88;
wire [0:0] new_89;
wire [0:0] new_90;
wire [0:0] new_91;
wire [0:0] new_92;
wire [0:0] new_93;
wire [0:0] new_94;
wire [0:0] new_95;
wire [0:0] new_96;
wire [0:0] new_97;
wire [0:0] new_98;
wire [0:0] new_99;
wire [0:0] new_100;
wire [0:0] new_101;
wire [0:0] new_102;
wire [0:0] new_103;
wire [0:0] new_104;
wire [0:0] new_106;
wire [0:0] new_107;
wire [0:0] new_108;
assign new_108 = i[5] ? 0 : 0;
assign new_107 = i[5] ? 0 : 0;
assign new_106 = i[9] ? 0 : 0;
assign new_104 = i[9] ? 0 : 0;
assign new_103 = i[8] ? 0 : 0;
assign new_102 = i[4] ? 0 : 0;
assign new_101 = i[5] ? 0 : 0;
assign new_100 = i[4] ? 0 : 0;
assign new_99 = i[4] ? 0 : 0;
assign new_98 = i[5] ? 0 : 0;
assign new_97 = i[5] ? 0 : 0;
assign new_96 = i[3] ? 0 : 0;
assign new_95 = i[4] ? 0 : 0;
assign new_94 = i[4] ? 0 : 0;
assign new_93 = i[10] ? 0 : 0;
assign new_92 = i[4] ? 0 : 0;
assign new_91 = i[1] ? 0 : 0;
assign new_90 = i[1] ? 0 : 0;
assign new_89 = i[10] ? 0 : 0;
assign new_88 = i[3] ? 0 : 0;
assign new_87 = i[9] ? 0 : 0;
assign new_85 = i[1] ? 0 : 0;
assign new_84 = i[1] ? 0 : 0;
assign new_82 = i[1] ? 0 : 0;
assign new_81 = i[8] ? 0 : 0;
assign new_80 = i[9] ? 0 : 0;
assign new_79 = i[3] ? 0 : 0;
assign new_77 = i[5] ? 0 : 0;
assign new_76 = i[9] ? 0 : 0;
assign new_75 = i[0] ? 0 : 0;
assign new_74 = i[9] ? 0 : 0;
assign new_73 = i[4] ? 0 : 0;
assign new_72 = i[4] ? 0 : 0;
assign new_71 = i[10] ? 0 : 0;
assign new_70 = i[2] ? 0 : 0;
assign new_69 = i[5] ? 0 : 0;
assign new_68 = i[1] ? 0 : 0;
assign new_67 = i[1] ? 0 : 0;
assign new_66 = i[9] ? 0 : 0;
assign new_65 = i[8] ? 0 : 0;
assign new_63 = i[3] ? 0 : 0;
assign new_61 = i[8] ? 0 : 0;
assign new_60 = i[8] ? 0 : 0;
assign new_59 = i[8] ? 0 : 0;
assign new_57 = i[42] ? 0 : 0;
assign new_55 = i[8] ? new_107 : new_108;
assign new_54 = i[5] ? 0 : new_106;
assign new_53 = i[5] ? new_103 : new_104;
assign new_52 = i[8] ? new_101 : new_102;
assign new_51 = i[3] ? new_99 : new_100;
assign new_50 = i[3] ? new_97 : new_98;
assign new_49 = i[0] ? new_95 : new_96;
assign new_48 = i[0] ? new_93 : new_94;
assign new_47 = i[3] ? new_91 : new_92;
assign new_46 = i[3] ? new_89 : new_90;
assign new_45 = i[1] ? new_87 : new_88;
assign new_44 = i[0] ? new_85 : 0;
assign new_43 = i[8] ? 0 : new_84;
assign new_42 = i[0] ? new_81 : new_82;
assign new_41 = i[1] ? new_79 : new_80;
assign new_40 = i[4] ? new_77 : 0;
assign new_39 = i[5] ? new_75 : new_76;
assign new_38 = i[8] ? new_73 : new_74;
assign new_37 = i[3] ? new_71 : new_72;
assign new_36 = i[4] ? new_69 : new_70;
assign new_34 = i[9] ? new_67 : new_68;
assign new_33 = i[1] ? new_65 : new_66;
assign new_32 = i[8] ? new_63 : 0;
assign new_31 = i[21] ? new_61 : 0;
assign new_30 = i[0] ? new_59 : new_60;
assign new_29 = i[44] ? new_57 : 0;
assign new_28 = i[0] ? new_55 : 0;
assign new_27 = i[0] ? new_53 : new_54;
assign new_26 = i[0] ? new_51 : new_52;
assign new_25 = i[8] ? new_49 : new_50;
assign new_24 = i[9] ? new_47 : new_48;
assign new_23 = i[5] ? new_45 : new_46;
assign new_22 = i[3] ? new_43 : new_44;
assign new_21 = i[4] ? new_41 : new_42;
assign new_20 = i[8] ? new_39 : new_40;
assign new_19 = i[0] ? new_37 : new_38;
assign new_18 = i[6] ? 0 : new_36;
assign new_17 = i[48] ? new_33 : new_34;
assign new_16 = i[37] ? new_31 : new_32;
assign new_15 = i[39] ? new_29 : new_30;
assign new_14 = i[4] ? new_27 : new_28;
assign new_13 = i[9] ? new_25 : new_26;
assign new_11 = i[8] ? new_23 : new_24;
assign new_10 = i[2] ? new_21 : new_22;
assign new_9 = i[1] ? new_19 : new_20;
assign new_8 = i[10] ? new_17 : new_18;
assign new_7 = i[1] ? new_15 : new_16;
assign new_6 = i[1] ? new_13 : new_14;
assign new_5 = i[2] ? new_11 : 0;
assign new_4 = i[49] ? new_9 : new_10;
assign new_3 = i[47] ? new_7 : new_8;
assign new_2 = i[48] ? new_5 : new_6;
assign new_1 = i[46] ? new_3 : new_4;
assign o = i[45] ? new_1 : new_2;


endmodule
