module class1_tree6(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_36;
wire [0:0] new_37;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_44;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_51;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_57;
wire [0:0] new_58;
wire [0:0] new_59;
wire [0:0] new_62;
wire [0:0] new_64;
wire [0:0] new_65;
assign new_65 = i[5] ? 0 : 0;
assign new_64 = i[5] ? 0 : 0;
assign new_62 = i[1] ? 0 : 0;
assign new_59 = i[1] ? 0 : 0;
assign new_58 = i[8] ? 0 : 0;
assign new_57 = i[1] ? 0 : 0;
assign new_55 = i[9] ? 0 : 0;
assign new_54 = i[9] ? 0 : 0;
assign new_53 = i[3] ? 0 : 0;
assign new_51 = i[3] ? 0 : 0;
assign new_47 = i[3] ? 0 : 0;
assign new_46 = i[0] ? 0 : 0;
assign new_45 = i[0] ? 0 : 0;
assign new_44 = i[8] ? 0 : 0;
assign new_43 = i[27] ? 0 : 0;
assign new_42 = i[46] ? 0 : 0;
assign new_41 = i[4] ? 0 : 0;
assign new_40 = i[4] ? 0 : 0;
assign new_39 = i[31] ? 0 : 0;
assign new_38 = i[4] ? new_65 : 0;
assign new_37 = i[1] ? 0 : new_64;
assign new_36 = i[4] ? 0 : new_62;
assign new_35 = i[5] ? new_59 : 0;
assign new_34 = i[4] ? new_57 : new_58;
assign new_33 = i[8] ? new_55 : 0;
assign new_31 = i[5] ? new_53 : new_54;
assign new_30 = i[5] ? new_51 : 0;
assign new_28 = i[8] ? 0 : 0;
assign new_27 = i[1] ? new_47 : 0;
assign new_26 = i[4] ? new_45 : new_46;
assign new_25 = i[10] ? new_43 : new_44;
assign new_24 = i[7] ? new_41 : new_42;
assign new_23 = i[40] ? new_39 : new_40;
assign new_21 = i[9] ? new_37 : new_38;
assign new_20 = i[9] ? new_35 : new_36;
assign new_19 = i[5] ? new_33 : new_34;
assign new_18 = i[1] ? new_31 : 0;
assign new_17 = i[8] ? 0 : new_30;
assign new_16 = i[4] ? new_27 : new_28;
assign new_14 = i[41] ? new_25 : new_26;
assign new_13 = i[10] ? new_23 : new_24;
assign new_12 = i[3] ? new_21 : 0;
assign new_10 = i[3] ? new_19 : new_20;
assign new_9 = i[4] ? new_17 : new_18;
assign new_8 = i[6] ? 0 : new_16;
assign new_7 = i[6] ? new_13 : new_14;
assign new_6 = i[48] ? 0 : new_12;
assign new_4 = i[0] ? new_9 : new_10;
assign new_3 = i[35] ? new_7 : new_8;
assign new_2 = i[8] ? 0 : new_6;
assign new_1 = i[17] ? new_3 : new_4;
assign o = i[42] ? new_1 : new_2;


endmodule
