module class1_tree1(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_36;
wire [0:0] new_37;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_44;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_49;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_52;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_56;
wire [0:0] new_57;
wire [0:0] new_59;
wire [0:0] new_60;
wire [0:0] new_61;
wire [0:0] new_63;
wire [0:0] new_64;
wire [0:0] new_65;
wire [0:0] new_66;
wire [0:0] new_67;
wire [0:0] new_68;
wire [0:0] new_69;
wire [0:0] new_70;
wire [0:0] new_72;
wire [0:0] new_73;
wire [0:0] new_74;
wire [0:0] new_75;
wire [0:0] new_77;
wire [0:0] new_78;
wire [0:0] new_80;
wire [0:0] new_81;
wire [0:0] new_84;
wire [0:0] new_86;
wire [0:0] new_87;
wire [0:0] new_88;
assign new_88 = i[6] ? 0 : 0;
assign new_87 = i[2] ? 0 : 0;
assign new_86 = i[9] ? 0 : 0;
assign new_84 = i[9] ? 0 : 0;
assign new_81 = i[2] ? 0 : 0;
assign new_80 = i[5] ? 0 : 0;
assign new_78 = i[1] ? 0 : 0;
assign new_77 = i[5] ? 0 : 0;
assign new_75 = i[4] ? 0 : 0;
assign new_74 = i[1] ? 0 : 0;
assign new_73 = i[36] ? 0 : 0;
assign new_72 = i[0] ? 0 : 0;
assign new_70 = i[0] ? 0 : 0;
assign new_69 = i[0] ? 0 : 0;
assign new_68 = i[0] ? 0 : 0;
assign new_67 = i[3] ? 0 : 0;
assign new_66 = i[2] ? 0 : 0;
assign new_65 = i[2] ? 0 : 0;
assign new_64 = i[6] ? 0 : 0;
assign new_63 = i[4] ? 0 : 0;
assign new_61 = i[4] ? 0 : 0;
assign new_60 = i[1] ? 0 : 0;
assign new_59 = i[5] ? 0 : 0;
assign new_57 = i[9] ? 0 : 0;
assign new_56 = i[4] ? 0 : 0;
assign new_55 = i[3] ? 0 : 0;
assign new_54 = i[4] ? 0 : 0;
assign new_53 = i[0] ? 0 : 0;
assign new_52 = i[1] ? 0 : 0;
assign new_51 = i[14] ? 0 : 0;
assign new_50 = i[1] ? 0 : 0;
assign new_49 = i[0] ? 0 : 0;
assign new_48 = i[3] ? new_87 : new_88;
assign new_47 = i[3] ? 0 : new_86;
assign new_46 = i[3] ? 0 : new_84;
assign new_45 = i[9] ? new_81 : 0;
assign new_44 = i[9] ? 0 : new_80;
assign new_43 = i[9] ? new_77 : new_78;
assign new_42 = i[9] ? new_75 : 0;
assign new_39 = i[26] ? new_73 : new_74;
assign new_38 = i[2] ? 0 : new_72;
assign new_37 = i[8] ? new_69 : new_70;
assign new_36 = i[2] ? new_67 : new_68;
assign new_35 = i[0] ? new_65 : new_66;
assign new_34 = i[5] ? new_63 : new_64;
assign new_33 = i[0] ? new_61 : 0;
assign new_32 = i[0] ? new_59 : new_60;
assign new_31 = i[4] ? new_57 : 0;
assign new_30 = i[48] ? new_55 : new_56;
assign new_29 = i[48] ? new_53 : new_54;
assign new_28 = i[31] ? new_51 : new_52;
assign new_27 = i[29] ? new_49 : new_50;
assign new_26 = i[8] ? new_47 : new_48;
assign new_25 = i[6] ? new_45 : new_46;
assign new_24 = i[3] ? new_43 : new_44;
assign new_22 = i[8] ? 0 : new_42;
assign new_21 = i[42] ? new_39 : 0;
assign new_20 = i[4] ? new_37 : new_38;
assign new_19 = i[8] ? new_35 : new_36;
assign new_18 = i[49] ? new_33 : new_34;
assign new_17 = i[49] ? new_31 : new_32;
assign new_16 = i[1] ? new_29 : new_30;
assign new_15 = i[49] ? new_27 : new_28;
assign new_14 = i[4] ? new_25 : new_26;
assign new_12 = i[0] ? 0 : new_24;
assign new_11 = i[47] ? new_21 : new_22;
assign new_9 = i[1] ? new_19 : new_20;
assign new_8 = i[8] ? new_17 : new_18;
assign new_7 = i[30] ? new_15 : new_16;
assign new_6 = i[0] ? 0 : new_14;
assign new_5 = i[45] ? new_11 : new_12;
assign new_4 = i[48] ? new_9 : 0;
assign new_3 = i[19] ? new_7 : new_8;
assign new_2 = i[46] ? new_5 : new_6;
assign new_1 = i[21] ? new_3 : new_4;
assign o = i[10] ? new_1 : new_2;


endmodule
