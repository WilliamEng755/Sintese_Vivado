module class0_tree3(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_3;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
assign new_32 = i[5] ? 0 : 0;
assign new_31 = i[4] ? 0 : 0;
assign new_30 = i[8] ? 0 : 0;
assign new_29 = i[1] ? 0 : 0;
assign new_28 = i[48] ? 0 : 0;
assign new_27 = i[9] ? 0 : 0;
assign new_26 = i[3] ? 0 : 0;
assign new_25 = i[3] ? 0 : 0;
assign new_24 = i[3] ? 0 : 0;
assign new_23 = i[8] ? 0 : 0;
assign new_22 = i[8] ? 0 : 0;
assign new_21 = i[0] ? 0 : 0;
assign new_20 = i[6] ? 0 : 0;
assign new_19 = i[14] ? 0 : 0;
assign new_18 = i[1] ? new_31 : new_32;
assign new_17 = i[4] ? new_29 : new_30;
assign new_16 = i[8] ? new_27 : new_28;
assign new_15 = i[9] ? new_25 : new_26;
assign new_14 = i[0] ? new_23 : new_24;
assign new_13 = i[1] ? new_21 : new_22;
assign new_11 = i[35] ? new_19 : new_20;
assign new_10 = i[3] ? new_17 : new_18;
assign new_9 = i[4] ? new_15 : new_16;
assign new_8 = i[10] ? new_13 : new_14;
assign new_7 = i[13] ? new_11 : 0;
assign new_6 = i[0] ? new_9 : new_10;
assign new_5 = i[45] ? new_7 : new_8;
assign new_3 = i[38] ? new_5 : new_6;
assign new_1 = i[12] ? new_3 : 0;
assign o = i[50] ? new_1 : 0;


endmodule
