module class1_tree0(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_36;
wire [0:0] new_37;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_49;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_56;
wire [0:0] new_58;
wire [0:0] new_59;
wire [0:0] new_60;
wire [0:0] new_61;
wire [0:0] new_62;
wire [0:0] new_63;
wire [0:0] new_64;
wire [0:0] new_65;
wire [0:0] new_66;
wire [0:0] new_67;
wire [0:0] new_68;
wire [0:0] new_69;
wire [0:0] new_70;
wire [0:0] new_71;
wire [0:0] new_72;
wire [0:0] new_74;
wire [0:0] new_75;
wire [0:0] new_78;
wire [0:0] new_79;
wire [0:0] new_80;
wire [0:0] new_81;
wire [0:0] new_83;
wire [0:0] new_84;
wire [0:0] new_85;
wire [0:0] new_86;
wire [0:0] new_87;
wire [0:0] new_88;
assign new_88 = i[3] ? 0 : 0;
assign new_87 = i[9] ? 0 : 0;
assign new_86 = i[4] ? 0 : 0;
assign new_85 = i[2] ? 0 : 0;
assign new_84 = i[6] ? 1 : 0;
assign new_83 = i[24] ? 0 : 0;
assign new_81 = i[3] ? 0 : 0;
assign new_80 = i[5] ? 0 : 0;
assign new_79 = i[5] ? 0 : 0;
assign new_78 = i[2] ? 0 : 0;
assign new_75 = i[4] ? 0 : 0;
assign new_74 = i[3] ? 0 : 0;
assign new_72 = i[5] ? 0 : 0;
assign new_71 = i[16] ? 0 : 0;
assign new_70 = i[4] ? 0 : 1;
assign new_69 = i[3] ? 0 : 0;
assign new_68 = i[3] ? 0 : 0;
assign new_67 = i[14] ? 0 : 0;
assign new_66 = i[1] ? 0 : 0;
assign new_65 = i[9] ? 0 : 1;
assign new_64 = i[1] ? 0 : 0;
assign new_63 = i[1] ? 0 : 0;
assign new_62 = i[10] ? 0 : 0;
assign new_61 = i[4] ? 0 : 0;
assign new_60 = i[0] ? 0 : 0;
assign new_59 = i[3] ? 0 : 0;
assign new_58 = i[0] ? 0 : 0;
assign new_56 = i[10] ? 1 : 0;
assign new_55 = i[49] ? 0 : 0;
assign new_54 = i[1] ? 0 : 0;
assign new_53 = i[30] ? 0 : 0;
assign new_51 = i[1] ? new_87 : new_88;
assign new_50 = i[6] ? new_85 : new_86;
assign new_49 = i[14] ? new_83 : new_84;
assign new_47 = i[4] ? new_81 : 0;
assign new_46 = i[3] ? new_79 : new_80;
assign new_45 = i[14] ? 0 : new_78;
assign new_41 = i[5] ? new_75 : 0;
assign new_40 = i[19] ? 0 : new_74;
assign new_39 = i[12] ? new_71 : new_72;
assign new_38 = i[5] ? new_69 : new_70;
assign new_37 = i[18] ? new_67 : new_68;
assign new_36 = i[5] ? new_65 : new_66;
assign new_35 = i[4] ? new_63 : new_64;
assign new_34 = i[1] ? new_61 : new_62;
assign new_32 = i[10] ? new_59 : new_60;
assign new_31 = i[1] ? 0 : new_58;
assign new_30 = i[1] ? new_55 : new_56;
assign new_29 = i[47] ? new_53 : new_54;
assign new_28 = i[4] ? new_51 : 0;
assign new_27 = i[18] ? new_49 : new_50;
assign new_26 = i[2] ? new_47 : 0;
assign new_25 = i[16] ? new_45 : new_46;
assign new_24 = i[5] ? 0 : 0;
assign new_23 = i[1] ? new_41 : 0;
assign new_22 = i[1] ? new_39 : new_40;
assign new_21 = i[19] ? new_37 : new_38;
assign new_18 = i[0] ? new_35 : new_36;
assign new_17 = i[0] ? 0 : new_34;
assign new_16 = i[8] ? new_31 : new_32;
assign new_15 = i[29] ? new_29 : new_30;
assign new_14 = i[16] ? new_27 : new_28;
assign new_13 = i[18] ? new_25 : new_26;
assign new_12 = i[9] ? new_23 : new_24;
assign new_11 = i[8] ? new_21 : new_22;
assign new_10 = i[4] ? 1 : 1;
assign new_8 = i[48] ? new_17 : new_18;
assign new_7 = i[46] ? new_15 : new_16;
assign new_6 = i[8] ? new_13 : new_14;
assign new_5 = i[23] ? new_11 : new_12;
assign new_4 = i[0] ? 1 : new_10;
assign new_3 = i[45] ? new_7 : new_8;
assign new_2 = i[0] ? new_5 : new_6;
assign new_1 = i[20] ? new_3 : new_4;
assign o = i[50] ? new_1 : new_2;


endmodule
