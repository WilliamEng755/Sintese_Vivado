module class5_tree0(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_15;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_26;
wire [0:0] new_27;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_36;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_44;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_49;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_52;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_56;
wire [0:0] new_57;
wire [0:0] new_58;
wire [0:0] new_59;
wire [0:0] new_61;
wire [0:0] new_63;
wire [0:0] new_64;
wire [0:0] new_65;
wire [0:0] new_66;
wire [0:0] new_67;
wire [0:0] new_69;
wire [0:0] new_70;
wire [0:0] new_71;
wire [0:0] new_72;
wire [0:0] new_73;
wire [0:0] new_74;
wire [0:0] new_75;
wire [0:0] new_77;
wire [0:0] new_78;
wire [0:0] new_79;
wire [0:0] new_80;
wire [0:0] new_81;
wire [0:0] new_82;
wire [0:0] new_83;
wire [0:0] new_84;
wire [0:0] new_85;
wire [0:0] new_86;
wire [0:0] new_87;
wire [0:0] new_88;
wire [0:0] new_89;
wire [0:0] new_90;
wire [0:0] new_91;
wire [0:0] new_93;
wire [0:0] new_94;
wire [0:0] new_96;
assign new_96 = i[5] ? 0 : 0;
assign new_94 = i[8] ? 0 : 0;
assign new_93 = i[4] ? 0 : 0;
assign new_91 = i[9] ? 0 : 1;
assign new_90 = i[3] ? 0 : 0;
assign new_89 = i[9] ? 0 : 0;
assign new_88 = i[0] ? 0 : 0;
assign new_87 = i[5] ? 0 : 0;
assign new_86 = i[1] ? 0 : 0;
assign new_85 = i[18] ? 0 : 0;
assign new_84 = i[6] ? 0 : 0;
assign new_83 = i[7] ? 0 : 0;
assign new_82 = i[3] ? 0 : 0;
assign new_81 = i[8] ? 0 : 0;
assign new_80 = i[9] ? 0 : 0;
assign new_79 = i[8] ? 0 : 1;
assign new_78 = i[8] ? 0 : 0;
assign new_77 = i[24] ? 0 : 0;
assign new_75 = i[4] ? 0 : 0;
assign new_74 = i[9] ? 0 : 0;
assign new_73 = i[9] ? 0 : 0;
assign new_72 = i[0] ? 0 : 0;
assign new_71 = i[0] ? 0 : 0;
assign new_70 = i[0] ? 0 : 0;
assign new_69 = i[9] ? 0 : 0;
assign new_67 = i[0] ? 0 : 0;
assign new_66 = i[9] ? 0 : 0;
assign new_65 = i[5] ? 0 : 0;
assign new_64 = i[9] ? 0 : 0;
assign new_63 = i[0] ? 0 : 0;
assign new_61 = i[5] ? 0 : 0;
assign new_59 = i[8] ? 0 : 0;
assign new_58 = i[5] ? 0 : 0;
assign new_57 = i[5] ? 0 : 0;
assign new_56 = i[5] ? 0 : 0;
assign new_55 = i[3] ? 0 : 0;
assign new_54 = i[1] ? 0 : 0;
assign new_53 = i[21] ? 0 : 0;
assign new_52 = i[9] ? 0 : new_96;
assign new_51 = i[3] ? new_93 : new_94;
assign new_50 = i[0] ? new_91 : 1;
assign new_49 = i[0] ? new_89 : new_90;
assign new_48 = i[9] ? new_87 : new_88;
assign new_47 = i[8] ? new_85 : new_86;
assign new_46 = i[8] ? new_83 : new_84;
assign new_45 = i[0] ? new_81 : new_82;
assign new_44 = i[1] ? new_79 : new_80;
assign new_43 = i[14] ? new_77 : new_78;
assign new_42 = i[0] ? new_75 : 0;
assign new_41 = i[0] ? new_73 : new_74;
assign new_40 = i[3] ? new_71 : new_72;
assign new_39 = i[3] ? new_69 : new_70;
assign new_38 = i[3] ? new_67 : 0;
assign new_36 = i[3] ? new_65 : new_66;
assign new_35 = i[2] ? new_63 : new_64;
assign new_34 = i[8] ? new_61 : 0;
assign new_32 = i[1] ? new_59 : 0;
assign new_31 = i[1] ? new_57 : new_58;
assign new_30 = i[1] ? new_55 : new_56;
assign new_29 = i[14] ? new_53 : new_54;
assign new_27 = i[0] ? new_51 : new_52;
assign new_26 = i[2] ? new_49 : new_50;
assign new_25 = i[2] ? new_47 : new_48;
assign new_24 = i[2] ? new_45 : new_46;
assign new_23 = i[19] ? new_43 : new_44;
assign new_22 = i[3] ? new_41 : new_42;
assign new_21 = i[4] ? new_39 : new_40;
assign new_20 = i[4] ? 0 : new_38;
assign new_19 = i[4] ? new_35 : new_36;
assign new_18 = i[0] ? 0 : new_34;
assign new_17 = i[0] ? new_31 : new_32;
assign new_15 = i[12] ? new_29 : new_30;
assign new_13 = i[2] ? new_27 : 0;
assign new_12 = i[15] ? new_25 : new_26;
assign new_11 = i[18] ? new_23 : new_24;
assign new_10 = i[1] ? new_21 : new_22;
assign new_9 = i[1] ? new_19 : new_20;
assign new_8 = i[3] ? new_17 : new_18;
assign new_7 = i[22] ? new_15 : 1;
assign new_6 = i[1] ? new_13 : 0;
assign new_5 = i[4] ? new_11 : new_12;
assign new_4 = i[8] ? new_9 : new_10;
assign new_3 = i[24] ? new_7 : new_8;
assign new_2 = i[13] ? new_5 : new_6;
assign new_1 = i[18] ? new_3 : new_4;
assign o = i[50] ? new_1 : new_2;


endmodule
