module class0_tree1(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_7;
wire [0:0] new_9;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_14;
wire [0:0] new_15;
wire [0:0] new_16;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_23;
wire [0:0] new_24;
wire [0:0] new_25;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_36;
wire [0:0] new_37;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_42;
assign new_42 = i[2] ? 0 : 0;
assign new_41 = i[0] ? 0 : 0;
assign new_40 = i[0] ? 0 : 0;
assign new_39 = i[6] ? 0 : 0;
assign new_37 = i[2] ? 0 : 0;
assign new_36 = i[9] ? 0 : 0;
assign new_35 = i[3] ? 0 : 0;
assign new_34 = i[1] ? 0 : 0;
assign new_33 = i[4] ? 0 : 0;
assign new_32 = i[3] ? 0 : 0;
assign new_31 = i[3] ? 0 : 0;
assign new_30 = i[8] ? 0 : 0;
assign new_29 = i[6] ? 0 : 0;
assign new_28 = i[0] ? 0 : 0;
assign new_27 = i[8] ? 0 : 0;
assign new_25 = i[46] ? 0 : 0;
assign new_24 = i[4] ? new_41 : new_42;
assign new_23 = i[4] ? new_39 : new_40;
assign new_21 = i[3] ? new_37 : 0;
assign new_20 = i[8] ? new_35 : new_36;
assign new_19 = i[8] ? new_33 : new_34;
assign new_18 = i[0] ? new_31 : new_32;
assign new_17 = i[48] ? new_29 : new_30;
assign new_16 = i[1] ? new_27 : new_28;
assign new_15 = i[28] ? new_25 : 1;
assign new_14 = i[1] ? new_23 : new_24;
assign new_13 = i[0] ? new_21 : 0;
assign new_12 = i[0] ? new_19 : new_20;
assign new_11 = i[1] ? new_17 : new_18;
assign new_9 = i[37] ? new_15 : new_16;
assign new_7 = i[8] ? new_13 : new_14;
assign new_6 = i[10] ? new_11 : new_12;
assign new_5 = i[12] ? new_9 : 0;
assign new_4 = i[48] ? new_7 : 1;
assign new_3 = i[31] ? new_5 : new_6;
assign new_1 = i[21] ? new_3 : new_4;
assign o = i[50] ? new_1 : 0;


endmodule
