module class5_tree2(input wire [50:0] i, output wire [0:0] o);

wire [0:0] new_1;
wire [0:0] new_2;
wire [0:0] new_3;
wire [0:0] new_4;
wire [0:0] new_5;
wire [0:0] new_6;
wire [0:0] new_8;
wire [0:0] new_9;
wire [0:0] new_10;
wire [0:0] new_11;
wire [0:0] new_12;
wire [0:0] new_13;
wire [0:0] new_15;
wire [0:0] new_17;
wire [0:0] new_18;
wire [0:0] new_19;
wire [0:0] new_20;
wire [0:0] new_21;
wire [0:0] new_22;
wire [0:0] new_23;
wire [0:0] new_25;
wire [0:0] new_27;
wire [0:0] new_28;
wire [0:0] new_29;
wire [0:0] new_30;
wire [0:0] new_31;
wire [0:0] new_32;
wire [0:0] new_33;
wire [0:0] new_34;
wire [0:0] new_35;
wire [0:0] new_37;
wire [0:0] new_38;
wire [0:0] new_39;
wire [0:0] new_40;
wire [0:0] new_41;
wire [0:0] new_42;
wire [0:0] new_43;
wire [0:0] new_44;
wire [0:0] new_45;
wire [0:0] new_46;
wire [0:0] new_47;
wire [0:0] new_48;
wire [0:0] new_50;
wire [0:0] new_51;
wire [0:0] new_52;
wire [0:0] new_53;
wire [0:0] new_54;
wire [0:0] new_55;
wire [0:0] new_56;
wire [0:0] new_57;
wire [0:0] new_58;
wire [0:0] new_59;
wire [0:0] new_60;
wire [0:0] new_61;
wire [0:0] new_63;
wire [0:0] new_64;
wire [0:0] new_65;
wire [0:0] new_66;
wire [0:0] new_67;
wire [0:0] new_68;
wire [0:0] new_69;
wire [0:0] new_70;
wire [0:0] new_71;
wire [0:0] new_72;
wire [0:0] new_73;
wire [0:0] new_74;
wire [0:0] new_75;
wire [0:0] new_76;
wire [0:0] new_77;
wire [0:0] new_78;
assign new_78 = i[4] ? 0 : 0;
assign new_77 = i[3] ? 0 : 0;
assign new_76 = i[5] ? 0 : 0;
assign new_75 = i[3] ? 0 : 0;
assign new_74 = i[4] ? 0 : 0;
assign new_73 = i[4] ? 0 : 0;
assign new_72 = i[5] ? 0 : 0;
assign new_71 = i[5] ? 0 : 0;
assign new_70 = i[3] ? 0 : 0;
assign new_69 = i[9] ? 0 : 0;
assign new_68 = i[0] ? 0 : 0;
assign new_67 = i[9] ? 0 : 0;
assign new_66 = i[5] ? 0 : 0;
assign new_65 = i[4] ? 0 : 0;
assign new_64 = i[8] ? 0 : 0;
assign new_63 = i[22] ? 0 : 0;
assign new_61 = i[5] ? 0 : 0;
assign new_60 = i[9] ? 0 : 0;
assign new_59 = i[5] ? 0 : 0;
assign new_58 = i[9] ? 0 : 0;
assign new_57 = i[9] ? 0 : 0;
assign new_56 = i[8] ? 0 : 0;
assign new_55 = i[4] ? 0 : 0;
assign new_54 = i[8] ? 0 : 0;
assign new_53 = i[6] ? 0 : 0;
assign new_52 = i[0] ? 0 : 0;
assign new_51 = i[6] ? 0 : 0;
assign new_50 = i[9] ? 0 : 0;
assign new_48 = i[0] ? 0 : 0;
assign new_47 = i[0] ? 0 : 0;
assign new_46 = i[1] ? 0 : 0;
assign new_45 = i[27] ? 0 : 0;
assign new_44 = i[9] ? new_77 : new_78;
assign new_43 = i[4] ? new_75 : new_76;
assign new_42 = i[2] ? new_73 : new_74;
assign new_41 = i[3] ? new_71 : new_72;
assign new_40 = i[0] ? new_69 : new_70;
assign new_39 = i[11] ? new_67 : new_68;
assign new_38 = i[8] ? new_65 : new_66;
assign new_37 = i[14] ? new_63 : new_64;
assign new_35 = i[4] ? new_61 : 0;
assign new_34 = i[0] ? new_59 : new_60;
assign new_33 = i[4] ? new_57 : new_58;
assign new_32 = i[0] ? new_55 : new_56;
assign new_31 = i[4] ? new_53 : new_54;
assign new_30 = i[2] ? new_51 : new_52;
assign new_29 = i[6] ? 0 : new_50;
assign new_28 = i[3] ? new_47 : new_48;
assign new_27 = i[12] ? new_45 : new_46;
assign new_25 = i[0] ? new_43 : new_44;
assign new_23 = i[0] ? new_41 : new_42;
assign new_22 = i[12] ? new_39 : new_40;
assign new_21 = i[11] ? new_37 : new_38;
assign new_20 = i[0] ? new_35 : 0;
assign new_19 = i[8] ? new_33 : new_34;
assign new_18 = i[9] ? new_31 : new_32;
assign new_17 = i[8] ? new_29 : new_30;
assign new_15 = i[24] ? new_27 : new_28;
assign new_13 = i[2] ? new_25 : 0;
assign new_12 = i[1] ? new_23 : 0;
assign new_11 = i[1] ? new_21 : new_22;
assign new_10 = i[3] ? new_19 : new_20;
assign new_9 = i[3] ? new_17 : new_18;
assign new_8 = i[23] ? new_15 : 1;
assign new_6 = i[1] ? new_13 : 0;
assign new_5 = i[15] ? new_11 : new_12;
assign new_4 = i[1] ? new_9 : new_10;
assign new_3 = i[49] ? 0 : new_8;
assign new_2 = i[13] ? new_5 : new_6;
assign new_1 = i[18] ? new_3 : new_4;
assign o = i[50] ? new_1 : new_2;


endmodule
